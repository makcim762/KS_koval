library verilog;
use verilog.vl_types.all;
entity ddnfv2 is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        q               : out    vl_logic
    );
end ddnfv2;
