module ddnfv2( 
  input x1, x2, x3, 
  output q 
); 
  assign q = (x1); 
endmodule


