module decoder4 (
    input  wire        en,       // Enable
    input  wire [3:0]  sel,      // Selector 0..15
    output reg  [15:0] out       // Output C0..C15
);

always @(*) begin
    if (en) begin
        case (sel)
            4'd0:  out = 16'b0000_0000_0000_0001; // C0 = 1
            4'd1:  out = 16'b0000_0000_0000_0010; // C1 = 1
            4'd2:  out = 16'b0000_0000_0000_0100; // C2 = 1
            4'd3:  out = 16'b0000_0000_0000_1000; // C3 = 1
            4'd4:  out = 16'b0000_0000_0001_0000; // C4 = 1
            4'd5:  out = 16'b0000_0000_0010_0000; // C5 = 1
            4'd6:  out = 16'b0000_0000_0100_0000; // C6 = 1
            4'd7:  out = 16'b0000_0000_1000_0000; // C7 = 1
            4'd8:  out = 16'b0000_0001_0000_0000; // C8 = 1
            4'd9:  out = 16'b0000_0010_0000_0000; // C9 = 1
            4'd10: out = 16'b0000_0100_0000_0000; // C10 = 1
            4'd11: out = 16'b0000_1000_0000_0000; // C11 = 1
            4'd12: out = 16'b0001_0000_0000_0000; // C12 = 1
            4'd13: out = 16'b0010_0000_0000_0000; // C13 = 1
            4'd14: out = 16'b0100_0000_0000_0000; // C14 = 1
            4'd15: out = 16'b1000_0000_0000_0000; // C15 = 1
            default: out = 16'b0000_0000_0000_0000;
        endcase
    end else begin
        out = 16'b0000_0000_0000_0000;
    end
end

endmodule
